package alu_uvm_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "alu_transaction.sv"
    `include "alu_driver.sv"
    `include "alu_monitor.sv"
    `include "alu_scoreboard.sv"
    `include "alu_agent.sv"
    `include "alu_env.sv"
    `include "alu_sequence.sv"
    `include "alu_random_test.sv"
endpackage